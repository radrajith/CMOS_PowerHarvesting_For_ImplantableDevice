** Profile: "SCHEMATIC1-sim"  [ C:\USERS\RADRA\BOX SYNC\SENIOR FALL 2016\ESE 440\Circuit simulation 1\laser sim1-PSpiceFiles\SCHEMATIC1\sim.sim ] 

** Creating circuit file "sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\radra\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V3 0 5 .1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
